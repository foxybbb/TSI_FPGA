--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   17:58:26 11/03/2022
-- Design Name:   
-- Module Name:   C:/Users/Ivan/Documents/FPGA/Pract_2/testdiv.vhd
-- Project Name:  Pract_2
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: frqDiv2
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY testdiv IS
END testdiv;
 
ARCHITECTURE behavior OF testdiv IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT frqDiv2
    PORT(
         D_IN : IN  std_logic;
         CLK_IN : IN  std_logic;
         CK_OUT : OUT  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal D_IN : std_logic := '0';
   signal CLK_IN : std_logic := '0';

 	--Outputs
   signal CK_OUT : std_logic;

   -- Clock period definitions
   constant CLK_IN_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: frqDiv2 PORT MAP (
          D_IN => D_IN,
          CLK_IN => CLK_IN,
          CK_OUT => CK_OUT
        );

   -- Clock process definitions
   CLK_IN_process :process
   begin
		CLK_IN <= '0';
		wait for CLK_IN_period/2;
		CLK_IN <= '1';
		wait for CLK_IN_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

      wait for CLK_IN_period*10;

      -- insert stimulus here 

      wait;
   end process;

END;
