
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity sgm is
    Port ( SeL : in  STD_LOGIC_VECTOR (3 downto 0);
			  ckIn: in STD_LOGIC;
			  ckEn: in STD_LOGIC;
           Sg : out  STD_LOGIC_VECTOR (6 downto 0));
end sgm;

architecture Structural of sgm is


   signal Sgm2 : std_logic_vector(13 downto 0);
begin

with SeL(3 downto 0) select
Sgm2(13 downto 0) <= "11111100110000" when "0000001",
                   "11111101101101" when "0000010",
                   "11111101111001" when "0000011",
                   "11111100110011" when "0000100",
                   "11111101011011" when "0000101",
                   "11111101011111" when "0000110",
                   "11111101110010" when "0000111",
                   "11111101111111" when "0001000",
                   "11111101111011" when "0001001",
                   "01100001111110" when "0001010",
                   "01100000110000" when "0001011",
                   "01100001101101" when "0001100",
                   "01100001111001" when "0001101",
                   "01100000110011" when "0001110",
                   "01100001011011" when "0001111",
                   "01100001011111" when "0010000",
                   "01100001110010" when "0010001",
                   "01100001111111" when "0010010",
                   "01100001111011" when "0010011",
                   "11011011111110" when "0010100",
                   "11011010110000" when "0010101",
                   "11011011101101" when "0010110",
                   "11011011111001" when "0010111",
                   "11011010110011" when "0011000",
                   "11011011011011" when "0011001",
                   "11011011011111" when "0011010",
                   "11011011110010" when "0011011",
                   "11011011111111" when "0011100",
                   "11011011111011" when "0011101",
                   "11110011111110" when "0011110",
                   "11110010110000" when "0011111",
                   "11110011101101" when "0100000",
                   "11110011111001" when "0100001",
                   "11110010110011" when "0100010",
                   "11110011011011" when "0100011",
                   "11110011011111" when "0100100",
                   "11110011110010" when "0100101",
                   "11110011111111" when "0100110",
                   "11110011111011" when "0100111",
                   "01100111111110" when "0101000",
                   "01100110110000" when "0101001",
                   "01100111101101" when "0101010",
                   "01100111111001" when "0101011",
                   "01100110110011" when "0101100",
                   "01100111011011" when "0101101",
                   "01100111011111" when "0101110",
                   "01100111110010" when "0101111",
                   "01100111111111" when "0110000",
                   "01100111111011" when "0110001",
                   "10110111111110" when "0110010",
                   "10110110110000" when "0110011",
                   "10110111101101" when "0110100",
                   "10110111111001" when "0110101",
                   "10110110110011" when "0110110",
                   "10110111011011" when "0110111",
                   "10110111011111" when "0111000",
                   "10110111110010" when "0111001",
                   "10110111111111" when "0111010",
                   "10110111111011" when "0111011",
                   "10111111111110" when "0111100",
                   "10111110110000" when "0111101",
                   "10111111101101" when "0111110",
                   "10111111111001" when "0111111",
                   "10111110110011" when "1000000",
                   "10111111011011" when "1000001",
                   "10111111011111" when "1000010",
                   "10111111110010" when "1000011",
                   "10111111111111" when "1000100",
                   "10111111111011" when "1000101",
                   "11100101111110" when "1000110",
                   "11100100110000" when "1000111",
                   "11100101101101" when "1001000",
                   "11100101111001" when "1001001",
                   "11100100110011" when "1001010",
                   "11100101011011" when "1001011",
                   "11100101011111" when "1001100",
                   "11100101110010" when "1001101",
                   "11100101111111" when "1001110",
                   "11100101111011" when "1001111",
                   "11111111111110" when "1010000",
                   "11111110110000" when "1010001",
                   "11111111101101" when "1010010",
                   "11111111111001" when "1010011",
                   "11111110110011" when "1010100",
                   "11111111011011" when "1010101",
                   "11111111011111" when "1010110",
                   "11111111110010" when "1010111",
                   "11111111111111" when "1011000",
                   "11111111111011" when "1011001",
                   "11110111111110" when "1011010",
                   "11110110110000" when "1011011",
                   "11110111101101" when "1011100",
                   "11110111111001" when "1011101",
                   "11110110110011" when "1011110",
                   "11110111011011" when "1011111",
                   "11110111011111" when "1100000",
                   "11110111110010" when "1100001",
                   "11110111111111" when "1100010",
                   "11110111111011" when "1100011",
                   "11111101111110" when others;

 Sgm0(6 downto 0) <= Sgm2(6 downto 0);
 Sgm1(13downto 0) <= Sgm2(13 downto 6);

 
process(ckIn)
begin
	if rising_edge(ckIn) then
		if ckEn = '1' then
		
		case (SeL) is 
      when "0001" =>Sg<="0110000";
      when "0010" =>Sg<="1101101";
      when "0011" =>Sg<="1111001";
      when "0100" =>Sg<="0110011";
      when "0101" =>Sg<="1011011";
      when "0110" =>Sg<="1011111";
      when "0111" =>Sg<="1110010";
      when "1000" =>Sg<="1111111";
      when "1001" =>Sg<="1111011";
      when "1010" =>Sg<="1110111";
      when "1011" =>Sg<="0011111";
      when "1100" =>Sg<="1001110";
      when "1101" =>Sg<="0111101";
      when "1110" =>Sg<="1001111";
      when "1111" =>Sg<="1000111";
      when others =>Sg<="1111110";
   end case;
		
		
		
		else
			
		end if;
	end if;
end process;



	 
end Structural;

